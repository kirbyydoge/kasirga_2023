`timescale 1ns/1ps
 
`include "sabitler.vh"

module crc16 (
    input clk_i,
    input rstn_i,
    input [7:0] byte_i,
    input  etkin_i,
    output [15:0] crc16_o
);
reg[15:0] tablo[255:0];

task tablo_init();
begin
   tablo[0] <= 16'h0000;
   tablo[1] <= 16'h1021;
   tablo[2] <= 16'h2042;
   tablo[3] <= 16'h3063;
   tablo[4] <= 16'h4084;
   tablo[5] <= 16'h50a5;
   tablo[6] <= 16'h60c6;
   tablo[7] <= 16'h70e7;
   tablo[8] <= 16'h8108;
   tablo[9] <= 16'h9129;
   tablo[10] <= 16'ha14a;
   tablo[11] <= 16'hb16b;
   tablo[12] <= 16'hc18c;
   tablo[13] <= 16'hd1ad;
   tablo[14] <= 16'he1ce;
   tablo[15] <= 16'hf1ef;
   tablo[16] <= 16'h1231;
   tablo[17] <= 16'h0210;
   tablo[18] <= 16'h3273;
   tablo[19] <= 16'h2252;
   tablo[20] <= 16'h52b5;
   tablo[21] <= 16'h4294;
   tablo[22] <= 16'h72f7;
   tablo[23] <= 16'h62d6;
   tablo[24] <= 16'h9339;
   tablo[25] <= 16'h8318;
   tablo[26] <= 16'hb37b;
   tablo[27] <= 16'ha35a;
   tablo[28] <= 16'hd3bd;
   tablo[29] <= 16'hc39c;
   tablo[30] <= 16'hf3ff;
   tablo[31] <= 16'he3de;
   tablo[32] <= 16'h2462;
   tablo[33] <= 16'h3443;
   tablo[34] <= 16'h0420;
   tablo[35] <= 16'h1401;
   tablo[36] <= 16'h64e6;
   tablo[37] <= 16'h74c7;
   tablo[38] <= 16'h44a4;
   tablo[39] <= 16'h5485;
   tablo[40] <= 16'ha56a;
   tablo[41] <= 16'hb54b;
   tablo[42] <= 16'h8528;
   tablo[43] <= 16'h9509;
   tablo[44] <= 16'he5ee;
   tablo[45] <= 16'hf5cf;
   tablo[46] <= 16'hc5ac;
   tablo[47] <= 16'hd58d;
   tablo[48] <= 16'h3653;
   tablo[49] <= 16'h2672;
   tablo[50] <= 16'h1611;
   tablo[51] <= 16'h0630;
   tablo[52] <= 16'h76d7;
   tablo[53] <= 16'h66f6;
   tablo[54] <= 16'h5695;
   tablo[55] <= 16'h46b4;
   tablo[56] <= 16'hb75b;
   tablo[57] <= 16'ha77a;
   tablo[58] <= 16'h9719;
   tablo[59] <= 16'h8738;
   tablo[60] <= 16'hf7df;
   tablo[61] <= 16'he7fe;
   tablo[62] <= 16'hd79d;
   tablo[63] <= 16'hc7bc;
   tablo[64] <= 16'h48c4;
   tablo[65] <= 16'h58e5;
   tablo[66] <= 16'h6886;
   tablo[67] <= 16'h78a7;
   tablo[68] <= 16'h0840;
   tablo[69] <= 16'h1861;
   tablo[70] <= 16'h2802;
   tablo[71] <= 16'h3823;
   tablo[72] <= 16'hc9cc;
   tablo[73] <= 16'hd9ed;
   tablo[74] <= 16'he98e;
   tablo[75] <= 16'hf9af;
   tablo[76] <= 16'h8948;
   tablo[77] <= 16'h9969;
   tablo[78] <= 16'ha90a;
   tablo[79] <= 16'hb92b;
   tablo[80] <= 16'h5af5;
   tablo[81] <= 16'h4ad4;
   tablo[82] <= 16'h7ab7;
   tablo[83] <= 16'h6a96;
   tablo[84] <= 16'h1a71;
   tablo[85] <= 16'h0a50;
   tablo[86] <= 16'h3a33;
   tablo[87] <= 16'h2a12;
   tablo[88] <= 16'hdbfd;
   tablo[89] <= 16'hcbdc;
   tablo[90] <= 16'hfbbf;
   tablo[91] <= 16'heb9e;
   tablo[92] <= 16'h9b79;
   tablo[93] <= 16'h8b58;
   tablo[94] <= 16'hbb3b;
   tablo[95] <= 16'hab1a;
   tablo[96] <= 16'h6ca6;
   tablo[97] <= 16'h7c87;
   tablo[98] <= 16'h4ce4;
   tablo[99] <= 16'h5cc5;
   tablo[100] <= 16'h2c22;
   tablo[101] <= 16'h3c03;
   tablo[102] <= 16'h0c60;
   tablo[103] <= 16'h1c41;
   tablo[104] <= 16'hedae;
   tablo[105] <= 16'hfd8f;
   tablo[106] <= 16'hcdec;
   tablo[107] <= 16'hddcd;
   tablo[108] <= 16'had2a;
   tablo[109] <= 16'hbd0b;
   tablo[110] <= 16'h8d68;
   tablo[111] <= 16'h9d49;
   tablo[112] <= 16'h7e97;
   tablo[113] <= 16'h6eb6;
   tablo[114] <= 16'h5ed5;
   tablo[115] <= 16'h4ef4;
   tablo[116] <= 16'h3e13;
   tablo[117] <= 16'h2e32;
   tablo[118] <= 16'h1e51;
   tablo[119] <= 16'h0e70;
   tablo[120] <= 16'hff9f;
   tablo[121] <= 16'hefbe;
   tablo[122] <= 16'hdfdd;
   tablo[123] <= 16'hcffc;
   tablo[124] <= 16'hbf1b;
   tablo[125] <= 16'haf3a;
   tablo[126] <= 16'h9f59;
   tablo[127] <= 16'h8f78;
   tablo[128] <= 16'h9188;
   tablo[129] <= 16'h81a9;
   tablo[130] <= 16'hb1ca;
   tablo[131] <= 16'ha1eb;
   tablo[132] <= 16'hd10c;
   tablo[133] <= 16'hc12d;
   tablo[134] <= 16'hf14e;
   tablo[135] <= 16'he16f;
   tablo[136] <= 16'h1080;
   tablo[137] <= 16'h00a1;
   tablo[138] <= 16'h30c2;
   tablo[139] <= 16'h20e3;
   tablo[140] <= 16'h5004;
   tablo[141] <= 16'h4025;
   tablo[142] <= 16'h7046;
   tablo[143] <= 16'h6067;
   tablo[144] <= 16'h83b9;
   tablo[145] <= 16'h9398;
   tablo[146] <= 16'ha3fb;
   tablo[147] <= 16'hb3da;
   tablo[148] <= 16'hc33d;
   tablo[149] <= 16'hd31c;
   tablo[150] <= 16'he37f;
   tablo[151] <= 16'hf35e;
   tablo[152] <= 16'h02b1;
   tablo[153] <= 16'h1290;
   tablo[154] <= 16'h22f3;
   tablo[155] <= 16'h32d2;
   tablo[156] <= 16'h4235;
   tablo[157] <= 16'h5214;
   tablo[158] <= 16'h6277;
   tablo[159] <= 16'h7256;
   tablo[160] <= 16'hb5ea;
   tablo[161] <= 16'ha5cb;
   tablo[162] <= 16'h95a8;
   tablo[163] <= 16'h8589;
   tablo[164] <= 16'hf56e;
   tablo[165] <= 16'he54f;
   tablo[166] <= 16'hd52c;
   tablo[167] <= 16'hc50d;
   tablo[168] <= 16'h34e2;
   tablo[169] <= 16'h24c3;
   tablo[170] <= 16'h14a0;
   tablo[171] <= 16'h0481;
   tablo[172] <= 16'h7466;
   tablo[173] <= 16'h6447;
   tablo[174] <= 16'h5424;
   tablo[175] <= 16'h4405;
   tablo[176] <= 16'ha7db;
   tablo[177] <= 16'hb7fa;
   tablo[178] <= 16'h8799;
   tablo[179] <= 16'h97b8;
   tablo[180] <= 16'he75f;
   tablo[181] <= 16'hf77e;
   tablo[182] <= 16'hc71d;
   tablo[183] <= 16'hd73c;
   tablo[184] <= 16'h26d3;
   tablo[185] <= 16'h36f2;
   tablo[186] <= 16'h0691;
   tablo[187] <= 16'h16b0;
   tablo[188] <= 16'h6657;
   tablo[189] <= 16'h7676;
   tablo[190] <= 16'h4615;
   tablo[191] <= 16'h5634;
   tablo[192] <= 16'hd94c;
   tablo[193] <= 16'hc96d;
   tablo[194] <= 16'hf90e;
   tablo[195] <= 16'he92f;
   tablo[196] <= 16'h99c8;
   tablo[197] <= 16'h89e9;
   tablo[198] <= 16'hb98a;
   tablo[199] <= 16'ha9ab;
   tablo[200] <= 16'h5844;
   tablo[201] <= 16'h4865;
   tablo[202] <= 16'h7806;
   tablo[203] <= 16'h6827;
   tablo[204] <= 16'h18c0;
   tablo[205] <= 16'h08e1;
   tablo[206] <= 16'h3882;
   tablo[207] <= 16'h28a3;
   tablo[208] <= 16'hcb7d;
   tablo[209] <= 16'hdb5c;
   tablo[210] <= 16'heb3f;
   tablo[211] <= 16'hfb1e;
   tablo[212] <= 16'h8bf9;
   tablo[213] <= 16'h9bd8;
   tablo[214] <= 16'habbb;
   tablo[215] <= 16'hbb9a;
   tablo[216] <= 16'h4a75;
   tablo[217] <= 16'h5a54;
   tablo[218] <= 16'h6a37;
   tablo[219] <= 16'h7a16;
   tablo[220] <= 16'h0af1;
   tablo[221] <= 16'h1ad0;
   tablo[222] <= 16'h2ab3;
   tablo[223] <= 16'h3a92;
   tablo[224] <= 16'hfd2e;
   tablo[225] <= 16'hed0f;
   tablo[226] <= 16'hdd6c;
   tablo[227] <= 16'hcd4d;
   tablo[228] <= 16'hbdaa;
   tablo[229] <= 16'had8b;
   tablo[230] <= 16'h9de8;
   tablo[231] <= 16'h8dc9;
   tablo[232] <= 16'h7c26;
   tablo[233] <= 16'h6c07;
   tablo[234] <= 16'h5c64;
   tablo[235] <= 16'h4c45;
   tablo[236] <= 16'h3ca2;
   tablo[237] <= 16'h2c83;
   tablo[238] <= 16'h1ce0;
   tablo[239] <= 16'h0cc1;
   tablo[240] <= 16'hef1f;
   tablo[241] <= 16'hff3e;
   tablo[242] <= 16'hcf5d;
   tablo[243] <= 16'hdf7c;
   tablo[244] <= 16'haf9b;
   tablo[245] <= 16'hbfba;
   tablo[246] <= 16'h8fd9;
   tablo[247] <= 16'h9ff8;
   tablo[248] <= 16'h6e17;
   tablo[249] <= 16'h7e36;
   tablo[250] <= 16'h4e55;
   tablo[251] <= 16'h5e74;
   tablo[252] <= 16'h2e93;
   tablo[253] <= 16'h3eb2;
   tablo[254] <= 16'h0ed1;
   tablo[255] <= 16'h1ef0;
end
endtask

reg[15:0] crc16_r,crc16_ns;
assign crc16_o = crc16_ns;
always@* begin
    crc16_ns = crc16_r;
    if(etkin_i) begin
        crc16_ns = {crc16_r<<8}^tablo[crc16_r[15:8]^byte_i];
    end
end

always@(posedge clk_i) begin
    if(!rstn_i) begin
        crc16_r <= 16'hffff;
        tablo_init();
    end else begin
        crc16_r <= crc16_ns;
    end
end

endmodule