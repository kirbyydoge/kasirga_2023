`define HUF_AC_0_0       16'b1010000000000000
`define HUF_AC_0_1       16'b0000000000000000
`define HUF_AC_0_2       16'b0100000000000000
`define HUF_AC_0_3       16'b1000000000000000
`define HUF_AC_0_4       16'b1011000000000000
`define HUF_AC_0_5       16'b1101000000000000
`define HUF_AC_0_6       16'b1111000000000000
`define HUF_AC_0_7       16'b1111100000000000
`define HUF_AC_0_8       16'b1111110110000000
`define HUF_AC_0_9       16'b1111111110000010
`define HUF_AC_0_10      16'b1111111110000011
`define HUF_AC_1_1       16'b1100000000000000
`define HUF_AC_1_2       16'b1101100000000000
`define HUF_AC_1_3       16'b1111001000000000
`define HUF_AC_1_4       16'b1111101100000000
`define HUF_AC_1_5       16'b1111111011000000
`define HUF_AC_1_6       16'b1111111110000100
`define HUF_AC_1_7       16'b1111111110000101
`define HUF_AC_1_8       16'b1111111110000110
`define HUF_AC_1_9       16'b1111111110000111
`define HUF_AC_1_10      16'b1111111110001000
`define HUF_AC_2_1       16'b1110000000000000
`define HUF_AC_2_2       16'b1111100100000000
`define HUF_AC_2_3       16'b1111110111000000
`define HUF_AC_2_4       16'b1111111101000000
`define HUF_AC_2_5       16'b1111111110001001
`define HUF_AC_2_6       16'b1111111110001010
`define HUF_AC_2_7       16'b1111111110001011
`define HUF_AC_2_8       16'b1111111110001100
`define HUF_AC_2_9       16'b1111111110001101
`define HUF_AC_2_10      16'b1111111110001110
`define HUF_AC_3_1       16'b1110100000000000
`define HUF_AC_3_2       16'b1111101110000000
`define HUF_AC_3_3       16'b1111111101010000
`define HUF_AC_3_4       16'b1111111110001111
`define HUF_AC_3_5       16'b1111111110010000
`define HUF_AC_3_6       16'b1111111110010001
`define HUF_AC_3_7       16'b1111111110010010
`define HUF_AC_3_8       16'b1111111110010011
`define HUF_AC_3_9       16'b1111111110010100
`define HUF_AC_3_10      16'b1111111110010101
`define HUF_AC_4_1       16'b1110110000000000
`define HUF_AC_4_2       16'b1111111000000000
`define HUF_AC_4_3       16'b1111111110010110
`define HUF_AC_4_4       16'b1111111110010111
`define HUF_AC_4_5       16'b1111111110011000
`define HUF_AC_4_6       16'b1111111110011001
`define HUF_AC_4_7       16'b1111111110011010
`define HUF_AC_4_8       16'b1111111110011011
`define HUF_AC_4_9       16'b1111111110011100
`define HUF_AC_4_10      16'b1111111110011101
`define HUF_AC_5_1       16'b1111010000000000
`define HUF_AC_5_2       16'b1111111011100000
`define HUF_AC_5_3       16'b1111111110011110
`define HUF_AC_5_4       16'b1111111110011111
`define HUF_AC_5_5       16'b1111111110100000
`define HUF_AC_5_6       16'b1111111110100001
`define HUF_AC_5_7       16'b1111111110100010
`define HUF_AC_5_8       16'b1111111110100011
`define HUF_AC_5_9       16'b1111111110100100
`define HUF_AC_5_10      16'b1111111110100101
`define HUF_AC_6_1       16'b1111011000000000
`define HUF_AC_6_2       16'b1111111101100000
`define HUF_AC_6_3       16'b1111111110100110
`define HUF_AC_6_4       16'b1111111110100111
`define HUF_AC_6_5       16'b1111111110101000
`define HUF_AC_6_6       16'b1111111110101001
`define HUF_AC_6_7       16'b1111111110101010
`define HUF_AC_6_8       16'b1111111110101011
`define HUF_AC_6_9       16'b1111111110101100
`define HUF_AC_6_10      16'b1111111110101101
`define HUF_AC_7_1       16'b1111101000000000
`define HUF_AC_7_2       16'b1111111101110000
`define HUF_AC_7_3       16'b1111111110101110
`define HUF_AC_7_4       16'b1111111110101111
`define HUF_AC_7_5       16'b1111111110110000
`define HUF_AC_7_6       16'b1111111110110001
`define HUF_AC_7_7       16'b1111111110110010 
`define HUF_AC_7_8       16'b1111111110110011
`define HUF_AC_7_9       16'b1111111110110100
`define HUF_AC_7_10      16'b1111111110110101
`define HUF_AC_8_1       16'b1111110000000000
`define HUF_AC_8_2       16'b1111111110000000
`define HUF_AC_8_3       16'b1111111110110110
`define HUF_AC_8_4       16'b1111111110110111
`define HUF_AC_8_5       16'b1111111110111000
`define HUF_AC_8_6       16'b1111111110111001
`define HUF_AC_8_7       16'b1111111110111010
`define HUF_AC_8_8       16'b1111111110111011
`define HUF_AC_8_9       16'b1111111110111100
`define HUF_AC_8_10      16'b1111111110111101
`define HUF_AC_9_1       16'b1111110010000000
`define HUF_AC_9_2       16'b1111111110111110
`define HUF_AC_9_3       16'b1111111110111111
`define HUF_AC_9_4       16'b1111111111000000
`define HUF_AC_9_5       16'b1111111111000001
`define HUF_AC_9_6       16'b1111111111000010
`define HUF_AC_9_7       16'b1111111111000011
`define HUF_AC_9_8       16'b1111111111000100
`define HUF_AC_9_9       16'b1111111111000101
`define HUF_AC_9_10      16'b1111111111000110
`define HUF_AC_10_1      16'b1111110100000000
`define HUF_AC_10_2      16'b1111111111000111
`define HUF_AC_10_3      16'b1111111111001000
`define HUF_AC_10_4      16'b1111111111001001
`define HUF_AC_10_5      16'b1111111111001010
`define HUF_AC_10_6      16'b1111111111001011
`define HUF_AC_10_7      16'b1111111111001100
`define HUF_AC_10_8      16'b1111111111001101
`define HUF_AC_10_9      16'b1111111111001110
`define HUF_AC_10_10     16'b1111111111001111
`define HUF_AC_11_1      16'b1111111001000000
`define HUF_AC_11_2      16'b1111111111010000
`define HUF_AC_11_3      16'b1111111111010001
`define HUF_AC_11_4      16'b1111111111010010
`define HUF_AC_11_5      16'b1111111111010011
`define HUF_AC_11_6      16'b1111111111010100
`define HUF_AC_11_7      16'b1111111111010101
`define HUF_AC_11_8      16'b1111111111010110
`define HUF_AC_11_9      16'b1111111111010111
`define HUF_AC_11_10     16'b1111111111011000
`define HUF_AC_12_1      16'b1111111010000000
`define HUF_AC_12_2      16'b1111111111011001
`define HUF_AC_12_3      16'b1111111111011010
`define HUF_AC_12_4      16'b1111111111011011
`define HUF_AC_12_5      16'b1111111111011100
`define HUF_AC_12_6      16'b1111111111011101
`define HUF_AC_12_7      16'b1111111111011110
`define HUF_AC_12_8      16'b1111111111011111
`define HUF_AC_12_9      16'b1111111111100000
`define HUF_AC_12_10     16'b1111111111100001
`define HUF_AC_13_1      16'b1111111100000000
`define HUF_AC_13_2      16'b1111111111100010
`define HUF_AC_13_3      16'b1111111111100011
`define HUF_AC_13_4      16'b1111111111100100
`define HUF_AC_13_5      16'b1111111111100101
`define HUF_AC_13_6      16'b1111111111100110
`define HUF_AC_13_7      16'b1111111111100111
`define HUF_AC_13_8      16'b1111111111101000
`define HUF_AC_13_9      16'b1111111111101001
`define HUF_AC_13_10     16'b1111111111101010
`define HUF_AC_14_1      16'b1111111111101011
`define HUF_AC_14_2      16'b1111111111101100
`define HUF_AC_14_3      16'b1111111111101101
`define HUF_AC_14_4      16'b1111111111101110
`define HUF_AC_14_5      16'b1111111111101111
`define HUF_AC_14_6      16'b1111111111110000
`define HUF_AC_14_7      16'b1111111111110001
`define HUF_AC_14_8      16'b1111111111110010
`define HUF_AC_14_9      16'b1111111111110011
`define HUF_AC_14_10     16'b1111111111110100
`define HUF_AC_15_1      16'b1111111111110101
`define HUF_AC_15_2      16'b1111111111110110
`define HUF_AC_15_3      16'b1111111111110111
`define HUF_AC_15_4      16'b1111111111111000
`define HUF_AC_15_5      16'b1111111111111001
`define HUF_AC_15_6      16'b1111111111111010
`define HUF_AC_15_7      16'b1111111111111011
`define HUF_AC_15_8      16'b1111111111111100
`define HUF_AC_15_9      16'b1111111111111101
`define HUF_AC_15_10     16'b1111111111111110
`define HUF_AC_15_0      16'b1111111100100000

`define EN_AC_0_0        16'b1111000000000000
`define EN_AC_0_1        16'b1100000000000000
`define EN_AC_0_2        16'b1100000000000000
`define EN_AC_0_3        16'b1110000000000000
`define EN_AC_0_4        16'b1111000000000000
`define EN_AC_0_5        16'b1111100000000000
`define EN_AC_0_6        16'b1111111000000000
`define EN_AC_0_7        16'b1111111100000000
`define EN_AC_0_8        16'b1111111111000000
`define EN_AC_0_9        16'b1111111111111111
`define EN_AC_0_10       16'b1111111111111111
`define EN_AC_1_1        16'b1111000000000000
`define EN_AC_1_2        16'b1111100000000000
`define EN_AC_1_3        16'b1111111000000000
`define EN_AC_1_4        16'b1111111110000000
`define EN_AC_1_5        16'b1111111111100000
`define EN_AC_1_6        16'b1111111111111111
`define EN_AC_1_7        16'b1111111111111111
`define EN_AC_1_8        16'b1111111111111111
`define EN_AC_1_9        16'b1111111111111111
`define EN_AC_1_10       16'b1111111111111111
`define EN_AC_2_1        16'b1111100000000000
`define EN_AC_2_2        16'b1111111100000000
`define EN_AC_2_3        16'b1111111111000000
`define EN_AC_2_4        16'b1111111111110000
`define EN_AC_2_5        16'b1111111111111111
`define EN_AC_2_6        16'b1111111111111111
`define EN_AC_2_7        16'b1111111111111111
`define EN_AC_2_8        16'b1111111111111111
`define EN_AC_2_9        16'b1111111111111111
`define EN_AC_2_10       16'b1111111111111111
`define EN_AC_3_1        16'b1111110000000000
`define EN_AC_3_2        16'b1111111110000000
`define EN_AC_3_3        16'b1111111111110000
`define EN_AC_3_4        16'b1111111111111111
`define EN_AC_3_5        16'b1111111111111111
`define EN_AC_3_6        16'b1111111111111111
`define EN_AC_3_7        16'b1111111111111111
`define EN_AC_3_8        16'b1111111111111111
`define EN_AC_3_9        16'b1111111111111111
`define EN_AC_3_10       16'b1111111111111111
`define EN_AC_4_1        16'b1111110000000000
`define EN_AC_4_2        16'b1111111111000000
`define EN_AC_4_3        16'b1111111111111111
`define EN_AC_4_4        16'b1111111111111111
`define EN_AC_4_5        16'b1111111111111111
`define EN_AC_4_6        16'b1111111111111111
`define EN_AC_4_7        16'b1111111111111111
`define EN_AC_4_8        16'b1111111111111111
`define EN_AC_4_9        16'b1111111111111111
`define EN_AC_4_10       16'b1111111111111111
`define EN_AC_5_1        16'b1111111000000000
`define EN_AC_5_2        16'b1111111111100000
`define EN_AC_5_3        16'b1111111111111111
`define EN_AC_5_4        16'b1111111111111111
`define EN_AC_5_5        16'b1111111111111111
`define EN_AC_5_6        16'b1111111111111111
`define EN_AC_5_7        16'b1111111111111111
`define EN_AC_5_8        16'b1111111111111111
`define EN_AC_5_9        16'b1111111111111111
`define EN_AC_5_10       16'b1111111111111111
`define EN_AC_6_1        16'b1111111000000000
`define EN_AC_6_2        16'b1111111111110000
`define EN_AC_6_3        16'b1111111111111111
`define EN_AC_6_4        16'b1111111111111111
`define EN_AC_6_5        16'b1111111111111111
`define EN_AC_6_6        16'b1111111111111111
`define EN_AC_6_7        16'b1111111111111111
`define EN_AC_6_8        16'b1111111111111111
`define EN_AC_6_9        16'b1111111111111111
`define EN_AC_6_10       16'b1111111111111111
`define EN_AC_7_1        16'b1111111100000000
`define EN_AC_7_2        16'b1111111111110000
`define EN_AC_7_3        16'b1111111111111111
`define EN_AC_7_4        16'b1111111111111111
`define EN_AC_7_5        16'b1111111111111111
`define EN_AC_7_6        16'b1111111111111111
`define EN_AC_7_7        16'b1111111111111111 
`define EN_AC_7_8        16'b1111111111111111
`define EN_AC_7_9        16'b1111111111111111
`define EN_AC_7_10       16'b1111111111111111
`define EN_AC_8_1        16'b1111111110000000
`define EN_AC_8_2        16'b1111111111111110
`define EN_AC_8_3        16'b1111111111111111
`define EN_AC_8_4        16'b1111111111111111
`define EN_AC_8_5        16'b1111111111111111
`define EN_AC_8_6        16'b1111111111111111
`define EN_AC_8_7        16'b1111111111111111
`define EN_AC_8_8        16'b1111111111111111
`define EN_AC_8_9        16'b1111111111111111
`define EN_AC_8_10       16'b1111111111111111
`define EN_AC_9_1        16'b1111111110000000
`define EN_AC_9_2        16'b1111111111111111
`define EN_AC_9_3        16'b1111111111111111
`define EN_AC_9_4        16'b1111111111111111
`define EN_AC_9_5        16'b1111111111111111
`define EN_AC_9_6        16'b1111111111111111
`define EN_AC_9_7        16'b1111111111111111
`define EN_AC_9_8        16'b1111111111111111
`define EN_AC_9_9        16'b1111111111111111
`define EN_AC_9_10       16'b1111111111111111
`define EN_AC_10_1       16'b1111111110000000
`define EN_AC_10_2       16'b1111111111111111
`define EN_AC_10_3       16'b1111111111111111
`define EN_AC_10_4       16'b1111111111111111
`define EN_AC_10_5       16'b1111111111111111
`define EN_AC_10_6       16'b1111111111111111
`define EN_AC_10_7       16'b1111111111111111
`define EN_AC_10_8       16'b1111111111111111
`define EN_AC_10_9       16'b1111111111111111
`define EN_AC_10_10      16'b1111111111111111
`define EN_AC_11_1       16'b1111111111000000
`define EN_AC_11_2       16'b1111111111111111
`define EN_AC_11_3       16'b1111111111111111
`define EN_AC_11_4       16'b1111111111111111
`define EN_AC_11_5       16'b1111111111111111
`define EN_AC_11_6       16'b1111111111111111
`define EN_AC_11_7       16'b1111111111111111
`define EN_AC_11_8       16'b1111111111111111
`define EN_AC_11_9       16'b1111111111111111
`define EN_AC_11_10      16'b1111111111111111
`define EN_AC_12_1       16'b1111111111000000
`define EN_AC_12_2       16'b1111111111111111
`define EN_AC_12_3       16'b1111111111111111
`define EN_AC_12_4       16'b1111111111111111
`define EN_AC_12_5       16'b1111111111111111
`define EN_AC_12_6       16'b1111111111111111
`define EN_AC_12_7       16'b1111111111111111
`define EN_AC_12_8       16'b1111111111111111
`define EN_AC_12_9       16'b1111111111111111
`define EN_AC_12_10      16'b1111111111111111
`define EN_AC_13_1       16'b1111111111100000
`define EN_AC_13_2       16'b1111111111111111
`define EN_AC_13_3       16'b1111111111111111
`define EN_AC_13_4       16'b1111111111111111
`define EN_AC_13_5       16'b1111111111111111
`define EN_AC_13_6       16'b1111111111111111
`define EN_AC_13_7       16'b1111111111111111
`define EN_AC_13_8       16'b1111111111111111
`define EN_AC_13_9       16'b1111111111111111
`define EN_AC_13_10      16'b1111111111111111
`define EN_AC_14_1       16'b1111111111111111
`define EN_AC_14_2       16'b1111111111111111
`define EN_AC_14_3       16'b1111111111111111
`define EN_AC_14_4       16'b1111111111111111
`define EN_AC_14_5       16'b1111111111111111
`define EN_AC_14_6       16'b1111111111111111
`define EN_AC_14_7       16'b1111111111111111
`define EN_AC_14_8       16'b1111111111111111
`define EN_AC_14_9       16'b1111111111111111
`define EN_AC_14_10      16'b1111111111111111
`define EN_AC_15_1       16'b1111111111111111
`define EN_AC_15_2       16'b1111111111111111
`define EN_AC_15_3       16'b1111111111111111
`define EN_AC_15_4       16'b1111111111111111
`define EN_AC_15_5       16'b1111111111111111
`define EN_AC_15_6       16'b1111111111111111
`define EN_AC_15_7       16'b1111111111111111
`define EN_AC_15_8       16'b1111111111111111
`define EN_AC_15_9       16'b1111111111111111
`define EN_AC_15_10      16'b1111111111111111
`define EN_AC_15_0       16'b1111111111100000

`define IDX_AC_0_0    'd0
`define IDX_AC_0_1    'd1
`define IDX_AC_0_2    'd2
`define IDX_AC_0_3    'd3
`define IDX_AC_0_4    'd4
`define IDX_AC_0_5    'd5
`define IDX_AC_0_6    'd6
`define IDX_AC_0_7    'd7
`define IDX_AC_0_8    'd8
`define IDX_AC_0_9    'd9
`define IDX_AC_0_10   'd10
`define IDX_AC_1_1    'd11
`define IDX_AC_1_2    'd12
`define IDX_AC_1_3    'd13
`define IDX_AC_1_4    'd14
`define IDX_AC_1_5    'd15
`define IDX_AC_1_6    'd16
`define IDX_AC_1_7    'd17
`define IDX_AC_1_8    'd18
`define IDX_AC_1_9    'd19
`define IDX_AC_1_10   'd20
`define IDX_AC_2_1    'd21
`define IDX_AC_2_2    'd22
`define IDX_AC_2_3    'd23
`define IDX_AC_2_4    'd24
`define IDX_AC_2_5    'd25
`define IDX_AC_2_6    'd26
`define IDX_AC_2_7    'd27
`define IDX_AC_2_8    'd28
`define IDX_AC_2_9    'd29
`define IDX_AC_2_10   'd30
`define IDX_AC_3_1    'd31
`define IDX_AC_3_2    'd32
`define IDX_AC_3_3    'd33
`define IDX_AC_3_4    'd34
`define IDX_AC_3_5    'd35
`define IDX_AC_3_6    'd36
`define IDX_AC_3_7    'd37
`define IDX_AC_3_8    'd38
`define IDX_AC_3_9    'd39
`define IDX_AC_3_10   'd40
`define IDX_AC_4_1    'd41
`define IDX_AC_4_2    'd42
`define IDX_AC_4_3    'd43
`define IDX_AC_4_4    'd44
`define IDX_AC_4_5    'd45
`define IDX_AC_4_6    'd46
`define IDX_AC_4_7    'd47
`define IDX_AC_4_8    'd48
`define IDX_AC_4_9    'd49
`define IDX_AC_4_10   'd50
`define IDX_AC_5_1    'd51
`define IDX_AC_5_2    'd52
`define IDX_AC_5_3    'd53
`define IDX_AC_5_4    'd54
`define IDX_AC_5_5    'd55
`define IDX_AC_5_6    'd56
`define IDX_AC_5_7    'd57
`define IDX_AC_5_8    'd58
`define IDX_AC_5_9    'd59
`define IDX_AC_5_10   'd60
`define IDX_AC_6_1    'd61
`define IDX_AC_6_2    'd62
`define IDX_AC_6_3    'd63
`define IDX_AC_6_4    'd64
`define IDX_AC_6_5    'd65
`define IDX_AC_6_6    'd66
`define IDX_AC_6_7    'd67
`define IDX_AC_6_8    'd68
`define IDX_AC_6_9    'd69
`define IDX_AC_6_10   'd70
`define IDX_AC_7_1    'd71
`define IDX_AC_7_2    'd72
`define IDX_AC_7_3    'd73
`define IDX_AC_7_4    'd74
`define IDX_AC_7_5    'd75
`define IDX_AC_7_6    'd76
`define IDX_AC_7_7    'd77
`define IDX_AC_7_8    'd78
`define IDX_AC_7_9    'd79
`define IDX_AC_7_10   'd80
`define IDX_AC_8_1    'd81
`define IDX_AC_8_2    'd82
`define IDX_AC_8_3    'd83
`define IDX_AC_8_4    'd84
`define IDX_AC_8_5    'd85
`define IDX_AC_8_6    'd86
`define IDX_AC_8_7    'd87
`define IDX_AC_8_8    'd88
`define IDX_AC_8_9    'd89
`define IDX_AC_8_10   'd90
`define IDX_AC_9_1    'd91
`define IDX_AC_9_2    'd92
`define IDX_AC_9_3    'd93
`define IDX_AC_9_4    'd94
`define IDX_AC_9_5    'd95
`define IDX_AC_9_6    'd96
`define IDX_AC_9_7    'd97
`define IDX_AC_9_8    'd98
`define IDX_AC_9_9    'd99
`define IDX_AC_9_10   'd100
`define IDX_AC_10_1   'd101
`define IDX_AC_10_2   'd102
`define IDX_AC_10_3   'd103
`define IDX_AC_10_4   'd104
`define IDX_AC_10_5   'd105
`define IDX_AC_10_6   'd106
`define IDX_AC_10_7   'd107
`define IDX_AC_10_8   'd108
`define IDX_AC_10_9   'd109
`define IDX_AC_10_10  'd110
`define IDX_AC_11_1   'd111
`define IDX_AC_11_2   'd112
`define IDX_AC_11_3   'd113
`define IDX_AC_11_4   'd114
`define IDX_AC_11_5   'd115
`define IDX_AC_11_6   'd116
`define IDX_AC_11_7   'd117
`define IDX_AC_11_8   'd118
`define IDX_AC_11_9   'd119
`define IDX_AC_11_10  'd120
`define IDX_AC_12_1   'd121
`define IDX_AC_12_2   'd122
`define IDX_AC_12_3   'd123
`define IDX_AC_12_4   'd124
`define IDX_AC_12_5   'd125
`define IDX_AC_12_6   'd126
`define IDX_AC_12_7   'd127
`define IDX_AC_12_8   'd128
`define IDX_AC_12_9   'd129
`define IDX_AC_12_10  'd130
`define IDX_AC_13_1   'd131
`define IDX_AC_13_2   'd132
`define IDX_AC_13_3   'd133
`define IDX_AC_13_4   'd134
`define IDX_AC_13_5   'd135
`define IDX_AC_13_6   'd136
`define IDX_AC_13_7   'd137
`define IDX_AC_13_8   'd138
`define IDX_AC_13_9   'd139
`define IDX_AC_13_10  'd140
`define IDX_AC_14_1   'd141
`define IDX_AC_14_2   'd142
`define IDX_AC_14_3   'd143
`define IDX_AC_14_4   'd144
`define IDX_AC_14_5   'd145
`define IDX_AC_14_6   'd146
`define IDX_AC_14_7   'd147
`define IDX_AC_14_8   'd148
`define IDX_AC_14_9   'd149
`define IDX_AC_14_10  'd150
`define IDX_AC_15_1   'd151
`define IDX_AC_15_2   'd152
`define IDX_AC_15_3   'd153
`define IDX_AC_15_4   'd154
`define IDX_AC_15_5   'd155
`define IDX_AC_15_6   'd156
`define IDX_AC_15_7   'd157
`define IDX_AC_15_8   'd158
`define IDX_AC_15_9   'd159
`define IDX_AC_15_10  'd160
`define IDX_AC_15_0   'd161

`define RUN_AC_0_0      4'd0   
`define RUN_AC_0_1      4'd0   
`define RUN_AC_0_2      4'd0   
`define RUN_AC_0_3      4'd0   
`define RUN_AC_0_4      4'd0   
`define RUN_AC_0_5      4'd0   
`define RUN_AC_0_6      4'd0   
`define RUN_AC_0_7      4'd0   
`define RUN_AC_0_8      4'd0   
`define RUN_AC_0_9      4'd0   
`define RUN_AC_0_10     4'd0  
`define RUN_AC_1_1      4'd1   
`define RUN_AC_1_2      4'd1   
`define RUN_AC_1_3      4'd1   
`define RUN_AC_1_4      4'd1   
`define RUN_AC_1_5      4'd1   
`define RUN_AC_1_6      4'd1   
`define RUN_AC_1_7      4'd1   
`define RUN_AC_1_8      4'd1   
`define RUN_AC_1_9      4'd1   
`define RUN_AC_1_10     4'd1  
`define RUN_AC_2_1      4'd2   
`define RUN_AC_2_2      4'd2   
`define RUN_AC_2_3      4'd2   
`define RUN_AC_2_4      4'd2   
`define RUN_AC_2_5      4'd2   
`define RUN_AC_2_6      4'd2   
`define RUN_AC_2_7      4'd2   
`define RUN_AC_2_8      4'd2   
`define RUN_AC_2_9      4'd2   
`define RUN_AC_2_10     4'd2  
`define RUN_AC_3_1      4'd3   
`define RUN_AC_3_2      4'd3   
`define RUN_AC_3_3      4'd3   
`define RUN_AC_3_4      4'd3   
`define RUN_AC_3_5      4'd3   
`define RUN_AC_3_6      4'd3   
`define RUN_AC_3_7      4'd3   
`define RUN_AC_3_8      4'd3   
`define RUN_AC_3_9      4'd3   
`define RUN_AC_3_10     4'd3  
`define RUN_AC_4_1      4'd4   
`define RUN_AC_4_2      4'd4   
`define RUN_AC_4_3      4'd4   
`define RUN_AC_4_4      4'd4   
`define RUN_AC_4_5      4'd4   
`define RUN_AC_4_6      4'd4   
`define RUN_AC_4_7      4'd4   
`define RUN_AC_4_8      4'd4   
`define RUN_AC_4_9      4'd4   
`define RUN_AC_4_10     4'd4  
`define RUN_AC_5_1      4'd5   
`define RUN_AC_5_2      4'd5   
`define RUN_AC_5_3      4'd5   
`define RUN_AC_5_4      4'd5   
`define RUN_AC_5_5      4'd5   
`define RUN_AC_5_6      4'd5   
`define RUN_AC_5_7      4'd5   
`define RUN_AC_5_8      4'd5   
`define RUN_AC_5_9      4'd5   
`define RUN_AC_5_10     4'd5  
`define RUN_AC_6_1      4'd6   
`define RUN_AC_6_2      4'd6   
`define RUN_AC_6_3      4'd6   
`define RUN_AC_6_4      4'd6   
`define RUN_AC_6_5      4'd6   
`define RUN_AC_6_6      4'd6   
`define RUN_AC_6_7      4'd6   
`define RUN_AC_6_8      4'd6   
`define RUN_AC_6_9      4'd6   
`define RUN_AC_6_10     4'd6  
`define RUN_AC_7_1      4'd7   
`define RUN_AC_7_2      4'd7   
`define RUN_AC_7_3      4'd7   
`define RUN_AC_7_4      4'd7   
`define RUN_AC_7_5      4'd7   
`define RUN_AC_7_6      4'd7   
`define RUN_AC_7_7      4'd7    
`define RUN_AC_7_8      4'd7   
`define RUN_AC_7_9      4'd7   
`define RUN_AC_7_10     4'd7  
`define RUN_AC_8_1      4'd8   
`define RUN_AC_8_2      4'd8   
`define RUN_AC_8_3      4'd8   
`define RUN_AC_8_4      4'd8   
`define RUN_AC_8_5      4'd8   
`define RUN_AC_8_6      4'd8   
`define RUN_AC_8_7      4'd8   
`define RUN_AC_8_8      4'd8   
`define RUN_AC_8_9      4'd8   
`define RUN_AC_8_10     4'd8  
`define RUN_AC_9_1      4'd9   
`define RUN_AC_9_2      4'd9   
`define RUN_AC_9_3      4'd9   
`define RUN_AC_9_4      4'd9   
`define RUN_AC_9_5      4'd9   
`define RUN_AC_9_6      4'd9   
`define RUN_AC_9_7      4'd9   
`define RUN_AC_9_8      4'd9   
`define RUN_AC_9_9      4'd9   
`define RUN_AC_9_10     4'd9  
`define RUN_AC_10_1     4'd10  
`define RUN_AC_10_2     4'd10  
`define RUN_AC_10_3     4'd10  
`define RUN_AC_10_4     4'd10  
`define RUN_AC_10_5     4'd10  
`define RUN_AC_10_6     4'd10  
`define RUN_AC_10_7     4'd10  
`define RUN_AC_10_8     4'd10  
`define RUN_AC_10_9     4'd10  
`define RUN_AC_10_10    4'd10 
`define RUN_AC_11_1     4'd11  
`define RUN_AC_11_2     4'd11  
`define RUN_AC_11_3     4'd11  
`define RUN_AC_11_4     4'd11  
`define RUN_AC_11_5     4'd11  
`define RUN_AC_11_6     4'd11  
`define RUN_AC_11_7     4'd11  
`define RUN_AC_11_8     4'd11  
`define RUN_AC_11_9     4'd11  
`define RUN_AC_11_10    4'd11 
`define RUN_AC_12_1     4'd12  
`define RUN_AC_12_2     4'd12  
`define RUN_AC_12_3     4'd12  
`define RUN_AC_12_4     4'd12  
`define RUN_AC_12_5     4'd12  
`define RUN_AC_12_6     4'd12  
`define RUN_AC_12_7     4'd12  
`define RUN_AC_12_8     4'd12  
`define RUN_AC_12_9     4'd12  
`define RUN_AC_12_10    4'd12 
`define RUN_AC_13_1     4'd13  
`define RUN_AC_13_2     4'd13  
`define RUN_AC_13_3     4'd13  
`define RUN_AC_13_4     4'd13  
`define RUN_AC_13_5     4'd13  
`define RUN_AC_13_6     4'd13  
`define RUN_AC_13_7     4'd13  
`define RUN_AC_13_8     4'd13  
`define RUN_AC_13_9     4'd13  
`define RUN_AC_13_10    4'd13 
`define RUN_AC_14_1     4'd14  
`define RUN_AC_14_2     4'd14  
`define RUN_AC_14_3     4'd14  
`define RUN_AC_14_4     4'd14  
`define RUN_AC_14_5     4'd14  
`define RUN_AC_14_6     4'd14  
`define RUN_AC_14_7     4'd14  
`define RUN_AC_14_8     4'd14  
`define RUN_AC_14_9     4'd14  
`define RUN_AC_14_10    4'd14 
`define RUN_AC_15_1     4'd15  
`define RUN_AC_15_2     4'd15  
`define RUN_AC_15_3     4'd15  
`define RUN_AC_15_4     4'd15  
`define RUN_AC_15_5     4'd15  
`define RUN_AC_15_6     4'd15  
`define RUN_AC_15_7     4'd15  
`define RUN_AC_15_8     4'd15  
`define RUN_AC_15_9     4'd15  
`define RUN_AC_15_10    4'd15 
`define RUN_AC_15_0     4'd15  

`define CAT_AC_0_0     4'd0   
`define CAT_AC_0_1     4'd1   
`define CAT_AC_0_2     4'd2   
`define CAT_AC_0_3     4'd3   
`define CAT_AC_0_4     4'd4   
`define CAT_AC_0_5     4'd5   
`define CAT_AC_0_6     4'd6   
`define CAT_AC_0_7     4'd7   
`define CAT_AC_0_8     4'd8   
`define CAT_AC_0_9     4'd9   
`define CAT_AC_0_10    4'd10  
`define CAT_AC_1_1     4'd1   
`define CAT_AC_1_2     4'd2   
`define CAT_AC_1_3     4'd3   
`define CAT_AC_1_4     4'd4   
`define CAT_AC_1_5     4'd5   
`define CAT_AC_1_6     4'd6   
`define CAT_AC_1_7     4'd7   
`define CAT_AC_1_8     4'd8   
`define CAT_AC_1_9     4'd9   
`define CAT_AC_1_10    4'd10  
`define CAT_AC_2_1     4'd1   
`define CAT_AC_2_2     4'd2   
`define CAT_AC_2_3     4'd3   
`define CAT_AC_2_4     4'd4   
`define CAT_AC_2_5     4'd5   
`define CAT_AC_2_6     4'd6   
`define CAT_AC_2_7     4'd7   
`define CAT_AC_2_8     4'd8   
`define CAT_AC_2_9     4'd9   
`define CAT_AC_2_10    4'd10  
`define CAT_AC_3_1     4'd1   
`define CAT_AC_3_2     4'd2   
`define CAT_AC_3_3     4'd3   
`define CAT_AC_3_4     4'd4   
`define CAT_AC_3_5     4'd5   
`define CAT_AC_3_6     4'd6   
`define CAT_AC_3_7     4'd7   
`define CAT_AC_3_8     4'd8   
`define CAT_AC_3_9     4'd9   
`define CAT_AC_3_10    4'd10  
`define CAT_AC_4_1     4'd1   
`define CAT_AC_4_2     4'd2   
`define CAT_AC_4_3     4'd3   
`define CAT_AC_4_4     4'd4   
`define CAT_AC_4_5     4'd5   
`define CAT_AC_4_6     4'd6   
`define CAT_AC_4_7     4'd7   
`define CAT_AC_4_8     4'd8   
`define CAT_AC_4_9     4'd9   
`define CAT_AC_4_10    4'd10  
`define CAT_AC_5_1     4'd1   
`define CAT_AC_5_2     4'd2   
`define CAT_AC_5_3     4'd3   
`define CAT_AC_5_4     4'd4   
`define CAT_AC_5_5     4'd5   
`define CAT_AC_5_6     4'd6   
`define CAT_AC_5_7     4'd7   
`define CAT_AC_5_8     4'd8   
`define CAT_AC_5_9     4'd9   
`define CAT_AC_5_10    4'd10  
`define CAT_AC_6_1     4'd1   
`define CAT_AC_6_2     4'd2   
`define CAT_AC_6_3     4'd3   
`define CAT_AC_6_4     4'd4   
`define CAT_AC_6_5     4'd5   
`define CAT_AC_6_6     4'd6   
`define CAT_AC_6_7     4'd7   
`define CAT_AC_6_8     4'd8   
`define CAT_AC_6_9     4'd9   
`define CAT_AC_6_10    4'd10  
`define CAT_AC_7_1     4'd1   
`define CAT_AC_7_2     4'd2   
`define CAT_AC_7_3     4'd3   
`define CAT_AC_7_4     4'd4   
`define CAT_AC_7_5     4'd5   
`define CAT_AC_7_6     4'd6   
`define CAT_AC_7_7     4'd7    
`define CAT_AC_7_8     4'd8   
`define CAT_AC_7_9     4'd9   
`define CAT_AC_7_10    4'd10  
`define CAT_AC_8_1     4'd1   
`define CAT_AC_8_2     4'd2   
`define CAT_AC_8_3     4'd3   
`define CAT_AC_8_4     4'd4   
`define CAT_AC_8_5     4'd5   
`define CAT_AC_8_6     4'd6   
`define CAT_AC_8_7     4'd7   
`define CAT_AC_8_8     4'd8   
`define CAT_AC_8_9     4'd9   
`define CAT_AC_8_10    4'd10  
`define CAT_AC_9_1     4'd1   
`define CAT_AC_9_2     4'd2   
`define CAT_AC_9_3     4'd3   
`define CAT_AC_9_4     4'd4   
`define CAT_AC_9_5     4'd5   
`define CAT_AC_9_6     4'd6   
`define CAT_AC_9_7     4'd7   
`define CAT_AC_9_8     4'd8   
`define CAT_AC_9_9     4'd9   
`define CAT_AC_9_10    4'd10  
`define CAT_AC_10_1    4'd1  
`define CAT_AC_10_2    4'd2  
`define CAT_AC_10_3    4'd3  
`define CAT_AC_10_4    4'd4  
`define CAT_AC_10_5    4'd5  
`define CAT_AC_10_6    4'd6  
`define CAT_AC_10_7    4'd7  
`define CAT_AC_10_8    4'd8  
`define CAT_AC_10_9    4'd9  
`define CAT_AC_10_10   4'd10 
`define CAT_AC_11_1    4'd1  
`define CAT_AC_11_2    4'd2  
`define CAT_AC_11_3    4'd3  
`define CAT_AC_11_4    4'd4  
`define CAT_AC_11_5    4'd5  
`define CAT_AC_11_6    4'd6  
`define CAT_AC_11_7    4'd7  
`define CAT_AC_11_8    4'd8  
`define CAT_AC_11_9    4'd9  
`define CAT_AC_11_10   4'd10 
`define CAT_AC_12_1    4'd1  
`define CAT_AC_12_2    4'd2  
`define CAT_AC_12_3    4'd3  
`define CAT_AC_12_4    4'd4  
`define CAT_AC_12_5    4'd5  
`define CAT_AC_12_6    4'd6  
`define CAT_AC_12_7    4'd7  
`define CAT_AC_12_8    4'd8  
`define CAT_AC_12_9    4'd9  
`define CAT_AC_12_10   4'd10 
`define CAT_AC_13_1    4'd1  
`define CAT_AC_13_2    4'd2  
`define CAT_AC_13_3    4'd3  
`define CAT_AC_13_4    4'd4  
`define CAT_AC_13_5    4'd5  
`define CAT_AC_13_6    4'd6  
`define CAT_AC_13_7    4'd7  
`define CAT_AC_13_8    4'd8  
`define CAT_AC_13_9    4'd9  
`define CAT_AC_13_10   4'd10 
`define CAT_AC_14_1    4'd1  
`define CAT_AC_14_2    4'd2  
`define CAT_AC_14_3    4'd3  
`define CAT_AC_14_4    4'd4  
`define CAT_AC_14_5    4'd5  
`define CAT_AC_14_6    4'd6  
`define CAT_AC_14_7    4'd7  
`define CAT_AC_14_8    4'd8  
`define CAT_AC_14_9    4'd9  
`define CAT_AC_14_10   4'd10 
`define CAT_AC_15_1    4'd1  
`define CAT_AC_15_2    4'd2  
`define CAT_AC_15_3    4'd3  
`define CAT_AC_15_4    4'd4  
`define CAT_AC_15_5    4'd5  
`define CAT_AC_15_6    4'd6  
`define CAT_AC_15_7    4'd7  
`define CAT_AC_15_8    4'd8  
`define CAT_AC_15_9    4'd9  
`define CAT_AC_15_10   4'd10 
`define CAT_AC_15_0    4'd0   

`define DQ_STEP_0      6'd1
`define DQ_STEP_1      6'd2
`define DQ_STEP_2      6'd9
`define DQ_STEP_3      6'd9