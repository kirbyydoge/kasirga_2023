`define N_ALPHA         2
`define N_COSINE        45

// `define ALPHA_ZERO      18'b000000000000000010
// `define ALPHA_NZ        18'b000000000000000100

// `define IDCT_COS_VAL0   18'b000000000000001000 
// `define IDCT_COS_VAL1   18'b000000000000000111 
// `define IDCT_COS_VAL2   18'b000000000000000110 
// `define IDCT_COS_VAL3   18'b000000000000000101 
// `define IDCT_COS_VAL4   18'b000000000000000100 
// `define IDCT_COS_VAL5   18'b000000000000000011 
// `define IDCT_COS_VAL6   18'b000000000000000001 
// `define IDCT_COS_VAL7   18'b111111111111111111 
// `define IDCT_COS_VAL8   18'b111111111111111011 
// `define IDCT_COS_VAL9   18'b111111111111111001 
// `define IDCT_COS_VAL10  18'b111111111111111100 
// `define IDCT_COS_VAL11  18'b111111111111111101 
// `define IDCT_COS_VAL12  18'b111111111111111010

// `define ALPHA_ZERO      24'b000000000000000010110101
// `define ALPHA_NZ        24'b000000000000000100000000

// `define IDCT_COS_VAL0   24'b000000000000001000000000
// `define IDCT_COS_VAL1   24'b000000000000000111110110
// `define IDCT_COS_VAL2   24'b000000000000000111011001
// `define IDCT_COS_VAL3   24'b000000000000000110101001
// `define IDCT_COS_VAL4   24'b000000000000000101101010
// `define IDCT_COS_VAL5   24'b000000000000000100011100
// `define IDCT_COS_VAL6   24'b000000000000000011000011
// `define IDCT_COS_VAL7   24'b000000000000000001100011
// `define IDCT_COS_VAL8   24'b111111111111111110011101
// `define IDCT_COS_VAL9   24'b111111111111111010010110
// `define IDCT_COS_VAL10  24'b111111111111111000001010
// `define IDCT_COS_VAL11  24'b111111111111111000100111
// `define IDCT_COS_VAL12  24'b111111111111111011100100
// `define IDCT_COS_VAL13  24'b111111111111111100111101
// `define IDCT_COS_VAL14  24'b111111111111111001010111

`define ALPHA_ZERO          32'b00000000000000000101101010000010
`define ALPHA_NZ            32'b00000000000000001000000000000000

`define IDCT_COS_VAL0       32'b00000000000000010000000000000000
`define IDCT_COS_VAL1       32'b00000000000000001111101100010100
`define IDCT_COS_VAL2       32'b00000000000000001110110010000011
`define IDCT_COS_VAL3       32'b00000000000000001101010011011011
`define IDCT_COS_VAL4       32'b00000000000000001011010100000100
`define IDCT_COS_VAL5       32'b00000000000000001000111000111001
`define IDCT_COS_VAL6       32'b00000000000000000110000111110111
`define IDCT_COS_VAL7       32'b00000000000000000011000111110001
`define IDCT_COS_VAL8       32'b11111111111111111100111000001111
`define IDCT_COS_VAL9       32'b11111111111111110100101011111100
`define IDCT_COS_VAL10      32'b11111111111111110000010011101100
`define IDCT_COS_VAL11      32'b11111111111111110001001101111101
`define IDCT_COS_VAL12      32'b11111111111111110111000111000111
`define IDCT_COS_VAL13      32'b11111111111111111001111000001001
`define IDCT_COS_VAL14      32'b11111111111111110010101100100101
