`define N_ALPHA         2
`define N_COSINE        45

`define ALPHA_ZERO      18'b000000000000000010
`define ALPHA_NZ        18'b000000000000000100

`define IDCT_COS_VAL0   18'b000000000000001000 
`define IDCT_COS_VAL1   18'b000000000000000111 
`define IDCT_COS_VAL2   18'b000000000000000110 
`define IDCT_COS_VAL3   18'b000000000000000101 
`define IDCT_COS_VAL4   18'b000000000000000100 
`define IDCT_COS_VAL5   18'b000000000000000011 
`define IDCT_COS_VAL6   18'b000000000000000001 
`define IDCT_COS_VAL7   18'b111111111111111111 
`define IDCT_COS_VAL8   18'b111111111111111011 
`define IDCT_COS_VAL9   18'b111111111111111001 
`define IDCT_COS_VAL10  18'b111111111111111100 
`define IDCT_COS_VAL11  18'b111111111111111101 
`define IDCT_COS_VAL12  18'b111111111111111010 
