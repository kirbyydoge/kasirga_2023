`timescale 1ns/1ps

`include "sabitler.vh"

module tb_top();

reg clk_i;
reg rstn_i;

reg  [7:0] rx_fifo_wr_data_w;
reg        rx_fifo_wr_en_w;
wire [7:0] rx_fifo_rd_data_w;
reg        rx_fifo_rd_en_w;
wire       rx_fifo_full_w;
wire       rx_fifo_empty_w;

fifo #(
   .DATA_WIDTH(8),
   .DATA_DEPTH(32)
) rx_buffer (
   .clk_i    ( clk_i ),         
   .rstn_i   ( rstn_i ),         
   .data_i   ( rx_fifo_wr_data_w ),         
   .wr_en_i  ( rx_fifo_wr_en_w ),         
   .data_o   ( rx_fifo_rd_data_w ),         
   .rd_en_i  ( rx_fifo_rd_en_w ),         
   .full_o   ( rx_fifo_full_w ),         
   .empty_o  ( rx_fifo_empty_w )         
);


wire[7:0] h_veri_i;
wire      h_gecerli_i;
wire     h_hazir_o;
wire[7:0] h_veri_o;
wire      h_gecerli_o;
wire      h_hazir_i;

assign h_veri_i = rx_fifo_rd_data_w;
assign h_gecerli_i = !rx_fifo_empty_w;
assign h_hazir_i = !tx_fifo_full_w;
assign rx_fifo_rd_en_w = h_hazir_o;

hizlandirici hz(
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .h_veri_i(h_veri_i),
    .h_gecerli_i(h_gecerli_i),
    .h_hazir_o(h_hazir_o),
    .h_veri_o(h_veri_o),
    .h_gecerli_o(h_gecerli_o),
    .h_hazir_i(h_hazir_i)
);

wire[7:0] rx_fifo_wr_data_w;
wire      rx_fifo_wr_en_w;
wire[7:0] tx_fifo_rd_data_w;
wire tx_fifo_rd_en_w;
wire tx_fifo_full_w;
wire tx_fifo_empty_w;

assign tx_fifo_wr_data_w = h_veri_o;
assign tx_fifo_wr_en_w = h_hazir_o;

fifo #(
   .DATA_WIDTH(8),
   .DATA_DEPTH(32)
) tx_buffer (
   .clk_i    ( clk_i ),         
   .rstn_i   ( rstn_i ),         
   .data_i   ( tx_fifo_wr_data_w ),         
   .wr_en_i  ( tx_fifo_wr_en_w ),         
   .data_o   ( tx_fifo_rd_data_w ),         
   .rd_en_i  ( tx_fifo_rd_en_w ),         
   .full_o   ( tx_fifo_full_w ),         
   .empty_o  ( tx_fifo_empty_w )         
);



always begin
    clk_i = 1'b1;
    #5;
    clk_i = 1'b0;
    #5;
end

localparam TEST_LEN = 34648;
localparam BYTE_LEN = TEST_LEN/8;
reg [TEST_LEN-1:0] temp_deger;
reg [7:0] bytes [0:BYTE_LEN-1];
localparam IMG_PATH ="D:/Teknofest_2023/kasirga-goruntu-2023/verify/tb_hd.txt";

integer step;

integer img_fd;
integer last_ctr;

always @(posedge clk_i) begin
    if (!rstn_i) begin
        last_ctr <= -1;
    end
    else if ( !tx_fifo_empty_w ) begin// && coz_hazir_i && last_ctr != denorm.dbg_ctr) begin
        $fwrite(img_fd, "%0d\n", tx_fifo_rd_data_w);
        $fflush(img_fd);
        tx_fifo_rd_en_w = 1;
    end else begin
        tx_fifo_rd_en_w = 0;
    end

end

integer i;
initial begin
    img_fd = $fopen(IMG_PATH, "w");
    step = 0;
    temp_deger = 34648'b1011101011001101_1010_0000_0001_0000_11101111101100000011110100000101000110000001111010000010100011000000111101000001010001100000011110100000101000110000001111010000010100011000000111101000001010001101101000111101000001010001100000011110100000111111001010100011000000111101000001010001100000011110100000101000110000001111010000010100011000000111101000001010001100000011110100000101000110000001111010000010100011000000111101000001010001100000011110100000101000110000001111010000010100011000000111101000001010001100000011110100000101000110000001111010000010100011000000111101000001010001100000011110100000101000110000001111010000010100011000000111101000001010001100000011110100000101000110000001111010000010100011000000111101000001010001100000011110100000101000110000001111010000010100011000000111101000001010001100000011110100000101000110000001111010000010100011000000111101000001010001100000011110100000101000110000001111010000010100011000000111101000001010001100000011110100000101000110000001111010000010100011000000111101000001010001100000011110100000101001011010001010001010010011001101000110011010001100110100011001101000110011010001100110100011001101000110011010001100110100100110011010001100110100011001101000110011010001100110100011001101000110011010001100110100011001101000110011010001100110100011001101000110011010001100110100011001101000110011010001100110100011001101000110011010001100110100101110011010001100110100011001101000110011010001100110100011001101000110011010001100110100100110011010001100110100011001101000110011010001100110100100110011010001100110100011001101000110011010010011001101000110011010001100110100011001101000110011010010011011101010001100110100011011101010001101110101000110111010100011011101010001101110101000110111010100011011101010001101110101000110111010100011011101010001101110101000110011010001100110100011001101001011100110100011001101000110011010001100110100101110011010001100110100011001101000110011010010111001101000110011010011011100110100011001101000110011010010011001101000110011010010011011101010001101110101001001101110101000110111010100100110111010100011011101010001101110101001001101110101000110111010100011011101010010011011101010001101110101000110111010100100110111010100011011101010001101110101000110111010100011011101010001101110101001011101110101000110111010100011011101010001101110101000110111010100101110111010100011011101010010111011101010001101110101000110111010100101110111010100011011101010010111011101010001101110101001011100110100011001101001101110111010100100110111010100100110111010100011011101010010011011101010010011011101010001101110101001001101110101001001101110101000110111110100100110111110100100110111110100011011111010010011011111010001101111101001001101111101000110111110100011011111010001101111101001001101111101000110111110100011011111010001101111101001011101111101000110111110100011011111010001101111101001011101111101000110111110100101110111110100011011111010010111011111010001101110101001011101110101001011101110101000110111010100101110111010100101110111010100011011101010010111011101010011001101110101001001101110101001001101110101001001101111101001001101111101001001101111101001000010111101001001101111101001001101111101001001101111101001001101111101000110111110100100110111110100100110111110100011011111010010011011111010001101111101000111100110010100100110111110100011011111010001101111101000110111110100011011111010001101111101000110111110100101110111110100011011111010010111011111010001101111101001011101111101001011101111101000110111110100101110111110100101110111110100101110111110100101110111110100101110111110100101110111010100101110111010100101110111010101000101101111101001000010111101001001101111101001000010111101001000010111101001101110111110100100001011110100100110111110100100110111110100100110111110100100001011110100100110111110100100110111110100011011111010010011011111010010011011111010001101111101000110111110100100110111110100011011111010001101111101000110111110100011011111010001101111101001011101111101000110111110100011011111010010111011111010010111011111010001101111101001011101111101001011101111101001010000111101001011101111101001011101111101001110110111110100101000011110100101000011110100101000011110100101000011110101000100010111101001000010111101001101001011110100100001011110100100001011110100110100101111010010011011111010011010010111101001001111001100101001001101111101001001101111101001001101111101001001101111101000110111110100100110111110100100110111110100011110011001010001101111101001001101111101000110111110100011011111010001101111101000110111110100011011111010010111011111010001101111101001011101111101000110111110100101110111110100101110111110100101111100110010100101000011110100101110111110100101000011110100101000011110100111000001111010010100001111010010100001111010011100000111101001010000111101010001000101111010011010010111101001000010111101001101001011110100100001011110100110100101111010011010010111101001000010111101001101001011110100100110111110100100110111110100100110111110100100110111110100011011111010010011110011001010011010011001001010010011110011011100010100101000100100110011010001101111110001010001111001100111101111010001111001100111101111010010111110011001010001101111101000110111110100111111110010001011101100001010011001110111010001000101101101100010000001101101011011001111001001001101001101110111110100011011111010010111011111010010111011111010000000111101001110000011110100101110111110100101110111110100101000011110100101000011110100111000001111010010100001111010011100000111101001010000111101001110000011110101000100010111101001101001011110100110100101111010011010010111101001000010111101001101001011110100110100101111010010011011111010010000101111010011010010111101001101110111110100110100101111010010011110011011010010111011111010011010010111001001111010010100101010101011001000011110011100011100010100111111011011111010100110100100110111001010101111011110100011011100000110000111010110101000100110110111000000111100000011100010100111001010010011100011101000011010011100001100100111101111010010111000001000111011110100110100100100100010100100111100111100111000000000110010011100000011101101100110100000010010110100101111100110010100101110111110100111000001101010010111011111010010111011111010010100001111010010100001111010011100000111101001010000111101001010000111101001110000011110100101000011110100111000001111010011100000111101010000100101111010010000101111010011010010111101001101001011110100100001011010100110100101101010011010010110101001101110111010100011011101010001100111001101000000010100100111101111010010111110010100000011111111000101010010000110001101000101111111100010101001101001010000001100011100000001101100010100111101011011011000001011110011111001100110010011010011110010010000101000110000000010010011010011000010100001011111111011101110010010011010100011001101101111001010000011100100111101001010010000101101101101111010110100101111110110110000101010001100000011011011111110010101010000101111011100101100111111111100010111111001010101000111101111100100001111110111011010011100000111100100010111111011110001101001011111001100001011011101111010100011001011111000001101001111010111011100011010011110001101110111011110100111100001101100010100101111100110010100011011111010010100001111010010100001111010011100000110101001110110111010100101110111110100101000011110100111000001111010011100000110101001010000111101001110000011110101000010010111101001000010111101001101001011110100100001011110100110111011101010010100000100100110101001000101100001011001111010100100000101100110010110111010010100001101011010000001000001100110010001110000000001010011010000001000011100111000010100111001111101111010100101010110110111010101111110100001111001101010000110111110100001010010110010100001111100110110010100010010010010011001111110111010100010011100011001111110101001111011010100110110110111100011100000100111100000111100110100000010010110001100011101001101101011100011101001111110001111011110100110101110101100001010100111100010010000111111100101010011000000010000000001100100000100100110101000000111101110110000101001110001100010100110100010111110011011111110000111100010100000110111010100110011100011100100100111000101001100110111100101101110101101001111000101101110010111111010000100010100110101111011001010011101011110010000001110001111011010100111010001110001110011001011110101111111010110100111000101000010110111010100100010100001011000110101000001111010110101001100001000111000110110000111000111000001101001111100101101100001011100110000100010010010011110010010010110001010001110110111000000001000010001010101001000011011011101110001111010111101011100110101010011010110011100111101110001010011110000011101111111010010100011011000110000111010110100110111001001000101001110000011010100111000001101010010111011111010010100001101010011100000110101001010000110101001110000011010100101000011010100111000001101010010100001101010100010001011010100100001011010100110100101101010000001100100100110101001000000101101001111000011001000100111010100110100100001101110010101000111010000110100011110011110110011011101000110001111111000010100001010101001011101101111100110110111001101010010001101011100110110100100010001110110100110010001001101110111101000000011100111111110010101001010011001011101111010111001100011100100111000111101010000011010100110110100111110011101101000011001110010011001110100111100111010001001101110101000001001111001000111101110001010101101111010100101011100100010111010000100011010110000110001011011000100010011100111111001100011110010010011010101010001010111100100000111000011001011000111100011111111011101101001010010101111100110011100011100000000010100111011111110110011101011011010010000011001011101110000000011111101001010100010100110101100011000001000000001100101010011000110001111011101100011111111010010101010010100101100110101101111000111110001101101011001111111011101010101110000001010101011000010111001101101010110001001110111011110011000100111111000011001101010111001000100001000111111001011000011110001001111101110010100111101110001010110100001001011101001110101111000010010101100110001100111111100101010110110010001010000010010001100111111011110111111110001101011001010101110111000101001110110001001011000000100100100011110110101010101000101001100110010100111000001000001101010010111011011001010111000110010101001101010001000110010010011110001000111111001100000011100011110101101010011110001110111010110010101110000010000000010001010011010111100101010111001111000010110101000111111001110001000001111000101001110111100111101101111010110100011110011100010011110110101001110000011011001101001110110111010100101000011010100111000001101010010100001101010010100001101010011100000110101001010000110101001110000011010100101000011010101000100010110101001001100100100110101001000100100011001001001111001101010110010001000000010000001110110000101010001010010000111011011110000001110010011010100000111100101010010010010100111000000000101010110001000111011001000001000001101110100100001110010011111010010101000111001011011101010000110001000111011000100000000011101111110110010101011111111010100111101101010100100101101111011001010011010111111011000000010111000011100101011000110011111111110010110011010111100000011111100011111010110101101010110000110110110110100010110110011011001101000101001010111010011011110100000111110011011000010111100000011110110110011110111001101011001111110101001110111010101100011101111010100010110111110000100010001011110011101110011011100011001111101101010101001101101011110110000010001001011100101101001111000100101000111111110111100001010101010010010011010111011011011101010110110110101001001000010111111110100000110000001111110101101001110101101111101010110010010011010010100001000111001011101000000011110100001111000001101001001011101110111011101110111100100100001010000011000110100111011011000111001001001111111000110101100111101100110011011001110111001100110011101101111101010011010011100101100111000001111111101111011001101010010001011011110011110010010011100001110111110000001111111011101111010110100111110010001111000101001101000010011001011000011000111100101100001110101000011000111111111000010101011000110100011110111111010001000011001000110101110011000010000110010101010101001110000100010000011000111110100111111101011010100111001110101110101011011100001100001000110101010011011000100000111110111010101001001110011100010101001100100101111110101000000110000010101110010001010010010010010010110001110011100011000010101010001100110101100111010111100111110110100110110011010100110010001010100011001100001111011010100101101101001101010101000100110000000000011101010001100100110101011010110111010001001110011100100101010101000101001111010100010110111011011101100001010000110100000100001001111110111011010100010001100000000111101101010100010011001010000100111011010101000110010111101001110100011110111010010001110101010001000001100101100110001110000000001010010101010010101011010010001110100100011011100001110010100000110010110001010100011100011000111110101101001010000110101001110000011010100111000001101010010100001101010010100001101010011100000110101001010000110101001100000001110010011010100110100011010111110110101010011001010110001010111111011101000110010011010010000100110010101100011110011110001010100100100011100001010011101010111011011001101010010110011010111001100001101101011000111100100000011001011000100011100001010001110101001101011000111100101101110011011100010111101100100110110111011101101101010000111101010000101101010110111011010010110011101101100101001000000001011100011011101111010010101101000110010001101011001110110110100010110011001011001110000101010100011111110000110001100111001001001101011100110111101010011110101010110011110011110010101110101101101010101110110001000010011100100011100011100100011111100011010110011010110100000101110011001000000010111100111100100000010000000111101010110100100011011000111111100111010100000011010001110110100010111100000110111011010000100111110110000001001101001100000011110110011010111111111100101101000110011011111010001011010000011011100110110111000001111110010100110010011111100000001010011100001011110111100000000001001011100001110101111101100110110010001010011101111001110101110001100011001000100100001011001011111101011100100010100110001111011101110011011000110000001100001011111011100000011100110101000100100011000100100111001001001110010011111011110101101100011010011000111010000101101101101001111010001101110101000101011101000011000011101001100100000111100101100101100101011000011100100011101010000011110010001010101001010011110110110101101100001001000110011010111001100100010001011001000001110010000111010100100000011011101111101010001111111010110101010011010110010110001101111001000110010110001110010001000011101101111010101100010011110000000001010101100010010100001011000110110000010110001100100101100000101111010101111111111011110001101001111100010101111011001000000011101100011101010101011010001111000111011111101010001010101010110111010100011100010110111111110011011000100100110000110111101101010101000101101001101001000000011110011010011111000111011101001100001110101101010111001000101001111100110001000110010101110111000010010001101010011100000101100011110111001111101000000001110111101010010101011011100000000101000000111010101101101110010000111100011001110001100010100111000101110000111000101010000001110100111101001010100100101100011011100100010110011101111001000111001110111100010111100110101000101110010000110010011001110001100100000100011000001111111100111010101101110111011101110111101001110010110000101111000111011000010110110100101010111011111110010010110011100100000011000111111000000011101011010110011110000110101001110000011010100111000001101010010100001101010011100000110101001010000110101001110000011010101001111000110100000000111001001101010010111011100001100011110100000101000111100110100000011101000001010011000011001011010011010011001101100000101010001100111000110010011100000011110111001101010110111001101101001100010100010110000011010111000100110011100101010011100111100111110111001111011000010101100000110111010101111101000101011010101010110010101110010000000010001110100010001011110111111110101001101011000110101110001101010110100110100111110010101000011011011010101111011000000011100000000010100100101101011101010111101110011011011010001011110010100010101010010010001011100111001000110111100011101001010011011001111101010111101110011001010001100001011101100100010000111111111010011001100011000001001111111000110101010001011001110110011101101100101100010010110001111101010011110011010011011100110100010100101000001110000011100110100111101010110110010011110100101010010001000110011110001101101100101000110110110111111010010101001010001001110001001001111100101100111000000000001001111010001100000001010011101111001011110000011111010100011101100010001010101100010000111011101000101110010101001001000001101011010110110100111110010010011010010101100000101000001001101011010011101111011111000011101100111101110011000100001001100100010100000111100011001001111001101011000111101101001011010010110101000100100100100010101111011101110001101000110000001000110000010000010000011100111100111001111010111101001010101111010111101101110001000111111101101000001000001001000010100101100110110000000101010111100110100110001110100110110011100001100011111100110000001110000010101110001110100111111000110100111011011111000000101100011110011001000111110110111001111010011001111011110101000101001101011001101011001000001101110010010101010001100101101101100110100011001111010010101011110110100111010111010101100111000101011011111111011001111011111110110100011010011001000000111110111101010110010000111100100000111100000011101001110111111010010100111111010100101011111110110101100111010101001000101011001010110111011010001010001101010011100100100101101100011001001111111000000010101010101010010010000111110101101010010111011110010011010010000100111001101001100101000110011010011100000011100110100111011001101001010000011010011100000011010010100001101010010100000110101011010110011010001110010011010011000111011100001011110001110111101001101010100001101001000011110001010110011101011101010111000011101011101010011100001010101001110010101100001001111001000111101010010011110101101010110011101011100110101111011111001011111110111001011101110101011011000001010000101000110001110010000001100011101110001010111001001010010010010001101001010110001011001110010010010010011010011001010001010001010001010001010001010010111011010010011110110101010010001010001100000000010100111010100100011100111011010101101001011000101001100111010011111011100001000110001111111011101011010101101010010110100100101100000101110000010000101011001110001000110111111011101010011111111010010101101111010110100111110110010110000001101000100101011110011001010101001011111111011101000000001111001011011111010010100111011010110111011111001011011110110111011101101111011000010110101001011011011000001000111100101101100001101100000101010010011110101000011011101101010101000101010011011000111010010110100011001101111101101011000011001100111110010000010101000010100001101110000001110111000001110001111111001010101010010111111111111011000100100101101001001101001001101111100011100101100100011000101110010011100100100100100000001100001010110101000101100001011100010110110101101100100110111101110111100011000010000011111101111000110000000110000101110011100111101110011110101001101001110000100101101100101011011101100010111010001000110101110011001010011111111000100110001111000000111111000111101011111110010110001010100000111111110001101111001001000110011100101100110110000001100100111101000000001100000000010100001100111000011100010101010101100100001110000011110100101001100000110000011010011100101000110000011010100101010110100111011100110100110100111001101001001010010100000110100111000000110100101000001101001110000001101001011100110100101110011010110100000000100110001010100011100100011111000111000000101001101100010100001001100100011011100111101001010110100011001100101100001110100111011010011110110101110001001000001100111001110010000101000111101011111111100111101001111110001101011100011111111111110111110101011101101101001011001111001111011101110010100111001001000000110111011111100011110110101011000111100100100100011010010001101101110011000111100110100110010100010100010100010100101000000110011110101111010010100111011001010100011101101010010011011100000001110100000101001001100100100111101111010011100101011111000111010111101001010100100010100100000111101001010010010010011111011100101010000110101001101000001001010000100001000000011000011111010001100001110101000101010110100000001001011011100010010001010110010100000101100110011001101101101010111000111101011010101100110011010011001001011011110000100110001001000011100100111111111100101101010111110011110010111001111101000001111011010101010111010110001110111010101110110100111111011101110110111010101010101001111010110010001100001100011001111111000100111101101111101001010100110111111111111100001001011000000010110111101110000100011110011110011010000001110100000001000001011001000000010010011100100011110100101011010000001100100010000000100111011000110001110110011111110000100000111101100001010010001010111000000001111110101101001110001000000111010110100111001000001110011110101101010010101101000000000111010111001101010000100110000011011011110111101001101001010111000101000110010010001010010100010010011110101101001110111000001000101001101001000110001010011011100110100111000000110100101110011010010100000110100111011001101001010000011010101110010010010111000111101000011010100010000011000101100110101011011010110100101110110001001100101011001010010111111010010101100101011110001010101101010000100010101110100101100101100010101101110011111110111010101101110010101100010000001000111011100111001001001001001111111010000010101110010011100111011100101011011010011011010001111111000100110111001111111000010101010010101000101000101001011100011110101001101001010000000000010011100000011001001001101010110100101110100111010111001011100000000100101010000100000001111111101111000111000101001011111101100001001010000111111001110111010100111110110000101001111000100010010000000011000110000001010011000110101101110100001010100100000011001000001111110101101010101000110010100101000110001000011000011100100010100001010110110110100111001101010010001111110010100001101010000110100010101101011110110101010000110110101101101000011001011110100100100100100000110000000011111111011101010111101110011010010011010011111011011101101011100110011001101001111101100110111001000100111000010001010011110100110011111010100110101011100001001100011011001111101101011011001100111011100111101010010010010010000101000111110100101010101000000000100010110010000101101000111100100101000010010011100011001111101001010100111010011001001000001110000000011100000011100111101001110110101001110000001101001111000011111100011000101001000011001000110010111100110100101100011101110110111000000111000001110010001010010101101011100000100111101011010011011111001101110011010011100000111000001101001011100010100101000110010001010011101110101101001100001010111000101001000000011010011100000011010011101100110100101110011010010100000110100111111100100100110101011101101100101000101100101110000010011010110101101001001011110001101011011010110010100111011110001111101010101100011001110001111101010011110000001111111001110101110001111101110101000010110100010110100101110001000100111111111100101101001001000010011100111110101110001111111111101011111001101011001010101111100011101101010110001010001111101111100011011100011111110001101010101001010010100000011001001000000101001110011000111100111000010111101001010100111101101111011010001101001001100001110110110000000101111111100111010101110110001001010101100001111001010100000000001101111010111000101001110001100100001001111010100100110100110100100100000110100110111100010100011100010100110101111000100100100100111010100011100111110101101010101101001001011010111011010001100100000110100110101010101000111100101101100000011110110101010001100101010001111010010101001111011001010110100011110111011101110010101100010100010010100101100010011010110111101101010011101101011000111001011111001011101101111000101001111011011110001001000101010100001011001001100010010111001111010011101111110110111011111110111101010101101111111111101100011000110011000001000101111001000000110111101001000110000001100100101011100011100100111110111001101000001100100001011010001100110001110001110001001011000100100001111010100111001110010110011011111010100110100110000010001111100011000101001101001100011011000000011000000110011100000110100111010001101010010101110011100111101001010011111010011010010010110000001110010000011110001111010010100111111011010000010001100100000011000101001001101100001001101001001101100001101000110001100010100111100000111110111101001110000011010100111000001101010010111001110011010010000100010100100101000110011010010111001101001010000011010101101001011100000000110101011110100000011011000010100011000101010110110110101101101111101101001101101000000101011100111011011000100010111110011001000110111101100001110110111111000110101100101011010110101000110110101110110101100010100010100001010000001010101010011100001010000001110100000000101011100111011101011001101100111001001011011101101000110010111000110010001101101110001100111101100011010110011001010011100101111000000001001111111001010100111000001001100000011001001101011010010101101110011100110110111010111110110111000101000011010100110110100100111001101000111001101000101001010001010010010010000011111001000011111101001010101011100000011000101001100110110000100101101101101000000110010011010110110110001000001111101100001101100010100100001010000111000100111100111010111011101001010011111111011101010111110100101010101011101001111100011000100110101110111111001100001000110011000111000011111100110111001111011100111101101111110101111111100101010101110111111111101111111011001010010111011001100110011100111011100110001001110010010010011010100000001011000011001101001000010011101110000110001010011110000000001111010000010100100001101000101001101001101001010101011000100010100111100001111010011111100100000110101000001001010000110011100111000000000110000001010010101010101110110001011100011001101001011100110100101000001101001110000001101001011101110101001011100110100010100010100101110011010100101010000100100101100001100110101101000010000100111111001011010101100011110011110010010100000010011001111000111101001010100110100011100011000001100010011000111000101011000001110101010110001100110011010000110010010001000101010010110001010100000101100101101011100101010011110101101010010100001010010001000110101001110001110101101010010110001001001111001100100100010101010010011100000000110101011110000010100001010101000010101010001100000000010100100001000101001100110001010010100000010100101110001010010111011011010001101101101000001010111001011001011110001111011010101010111000100010001011001101101101000111101011010101111010110101100011010110110110100101100010100100001100011000100110100100001011011001111100101111110101000101010011111010100101011100011111011010110110011100100000110001110001110010101111100011011100000101001001011000000000011110100110011010011001000011000110011011010110110111000100010011000100011011110111001110111001101110011111110010000101001000110101010001100100010100100000101010010001010011010010100100011001000101001001010001110000011010010000100010100100111010010100101110011010010111001101001000010011010010011001101001010000011010011100000011010010111001101001011100110100101110011010001100110100010101001101000111110101000101010111100101011011000010010100100111100110011000111011110101011110100000100111000011010001111000000101010001100010011110110110101100001001010001011101010111010000110111001010010110000010011111010011001111011110101010110100101110100001111010011011011111101011001101001101111100110101101110001101110000110110001110100001110111000000111001111111101001010110001101011101111010001111111001001001111100101001001011101010000001100110010100111101001100100111111110101000101010101110011011000110111001101101001100001111001011000010011101101111011001100001110010000011111110001101001111000111001111001000111011110100110101000010011100100101010110111001001111101011010011101101101111000110011010001101101000001101001011101101101001011101101101000110000000001110101101000000000011110010100100000010000110001101110111011011101101101101010100100110101001111000011011010001101000000000110011010111001100101010010000100000111101010001100011011100111111110100000000111011010101000101001011001000001101111111100101110000010001101111100101101111111000011110101011101101111101011111010010100101010110110110111100101100011011111001100110000110111011111111100111100110101001111000111111000100111101111010011001001001111110111100011011001001001111001101001001101110011001010000000001100111001101010010000011000011000011100000110100100001010111000101001000001010100100000001101001000010001010011000010010010001010010100001101010010110100100110001010010100010100000100010100110111000101000000101001110000001101001011100110100101110011010001100110100101110011010010111001101010110000101001000010110101001000011001011100100011000101010001101111001001010100100100000101110001101100001111010110100110110111000011101001011101110001101111000001001000011111100101011111101000011111010000111101100011010110000100101100110101110001011000110011100101010101100100011010001101100101001110000010001100111100011111100101111010010101001110101110101000011110011010110000111110110101000100101100111000111111111001011010001011110101111111000111110101101010110101000101011101110011001010010010110101101111001100001001000101001000111001000111010111111100110000011010010001111101100001010100001100111010100110000101100011110101110110100011001010111111100101110110101001100010110001111011100011100101011001011000110110000111101001100111000001111111010110101001010001000001001011111111110011110011001111111000011100110100101111110110001110011111101010001000010111110001111010111000101000000101101110010101111001011110010110000101001111011001101001001110011111110100110011010010001100110100000000110000101100011011101111001111001001111010001000101110000101111111001111101011010010001100001001111000110001101110001100101100000100001111101000000000010001100111111111000110101000110110101111101001000101010111000001101110101001011001001111011000000111000000101001011000011011010010111011101110010010001001001100111111011001111000101111111011111011111101011111110000111011100110101011010100100100100101101011011010001000011000111011011000000100100100111111011110011100111101010110111110101001101010100010110100100001011000110100011001101000111010110100111001010011100011101110011010011101100111001101000101001010001010011110101111001101001000110010010101000111101101101001011010010111000101000101001110101001000010001010011011010001010010100000110100101101000101001011010010110100111111001001001001101001111110111011000000101010000101101001001100100110101000110011001010010000011010011100101100100110011010011001011100101011000111011100001010000001001000101110010010001110000000110000111010100010101010001011110110010011101011110011000100110111100110000000011110100111000001000111111000010101000110000010010101011011001111001010101110001110111000111000001101010011111111011011101001111101101110110101110111110111100011110100011100011001111111010110100101010110111001100001111010101100101011001010011111011011100110101001000001001111000001110110011001110001111110010101001010011001110100110001100000001110111001000111101001100111000101001101000100101010100000111111001001000101100100111110111111001101010110011000111011001010111110101110000001100111000011010001101001111010101100011101101000101010010101001101001001101101010101001000111100111110111010001001001111011111011000001111111010100110101011000111100110011010011111011001001011111111010001111000101101111011100011111110001101111110010011111110000101010100011011100010111100100100100110011000111001001001110000011010101011111101011010011100001010010111000101001011010001010010100000110100111000000110100101000101001110010100111000101010010011011100000010001110011010011000110001000110011010011011100110100101110011010001010001010000011010011010011010010010100101101001010000011010010110100010100101101010010000100100001010001010100001011001111100110100110000100110100110010100101000001101001011100110100110111001001000001101001000111011000001111110000111000000011100011110111111010111111100111010100011000101101111011011100100111001011001101001010101111101101110001010011110001011011110110110111111111001111010101111111111110111110011010100100010110110111101100110001111111000101001000110111111001000010101001101000111111101100010010011101011000010010110111111110111100110001101010011000011010100000100100010000110001011011110000101000100111101110000101111001111111001110101010111100101101110111001111001010011100101100110001101010000100101110011111010111001001101001100111001001001111001101001011100010100101000000101001110000000101001011100010100011000101000110001010001100010100101101001011010010111001101001010000011010010000110100100101001010000011010010111001101001011100110100010100011000101001101001000101000101001011010001010010110100010100110101100110001001101001101101001001100011001101001000011010000001010010110100110000110100110101101110011010010011100100011101111010010111001111101100001010001101110111111110110010001010010111011101111111101100100010100101110111100111101100000000001010010000111001001111010100110100011000101001011100010100011000101001010001010011100001010010110100010100010100010100010100010100101101001010001010001010001010010010100101101001011010001010001100110100011001101000101000101000101000101001011010100011101000101001001010010000110100000010100101001111000000101001100001101001101101001001100010100101110001010001010001100010100111011000101001011100010100101110001010001100010100011000101000101001011010010110100010100010100010100100101001011010010110100010100101101000110011010001010001010001010010110100100101000101001011010001010001010001010001010011001010001010010000110100100101001110000000101001101011000110100110111000101001001100010100011000101001011100010100011000101001011100010100101110001010010110100010100010100010100010100010100010100101101000101000101000110001010010110100010100010100010100010100010100010100101101001011010000011010010010100010100101101000101000101000101001101110001010010000100110100110110100111000000010100000100110100110110100100110001010001100010100101000000101001011010010010100101101001011010001010010010100010100101101000101000101000101001011010001010001010001010001010001010010110100010100010100100101000101000101001011100110100101101001001010001010001010010110100010100010100000000;
    for (i = 0; i < BYTE_LEN; i = i + 1) begin
        bytes[i] = temp_deger[TEST_LEN - 1 - 8 * i -: 8];
    end
    rstn_i = 1'b0;
    rx_fifo_wr_en_w = 0;
    repeat(20) @(posedge clk_i);
    rstn_i = 1'b1;

    for (i = 0; i < BYTE_LEN;) begin
        rx_fifo_wr_data_w = bytes[i];
        rx_fifo_wr_en_w = 1;
        @(posedge clk_i); #2;
        if (!rx_fifo_full_w && !tx_fifo_full_w) begin
            i = i + 1;
        end
    end
    rx_fifo_wr_en_w = 1'b0;
end

endmodule