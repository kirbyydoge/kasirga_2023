`timescale 1ns/1ps

`include "sabitler.vh"

module tb_hd();

localparam TEST_AC_0_0   =  4'b1010;
localparam TEST_AC_0_1   =  2'b00;
localparam TEST_AC_0_2   =  2'b01;
localparam TEST_AC_0_3   =  3'b100;
localparam TEST_AC_0_4   =  4'b1011;
localparam TEST_AC_0_5   =  5'b11010;
localparam TEST_AC_0_6   =  7'b1111000;
localparam TEST_AC_0_7   =  8'b11111000;
localparam TEST_AC_0_8   = 10'b1111110110;
localparam TEST_AC_0_9   = 16'b1111111110000010;
localparam TEST_AC_0_10  = 16'b1111111110000011;

reg                       clk_i;
reg                       rstn_i;
reg     [`WB_BIT-1:0]     m_veri_i;
reg                       m_gecerli_i;
wire                      m_hazir_o;
wire    [10:0]            dc_data_o;
wire                      dc_valid_o;
reg                       dc_ready_i;
wire    [`RUN_BIT-1:0]    nd_run_o;
wire    [`HDATA_BIT-1:0]  nd_data_o;
wire    [`CAT_BIT-1:0]    nd_cat_o;
wire                      nd_gecerli_o;
wire                      nd_hazir_i;
wire                      nd_blk_son_o;

wire  [`HDATA_BIT-1:0]    ct_veri_o;
wire  [`BLOCK_BIT-1:0]    ct_row_o;
wire  [`BLOCK_BIT-1:0]    ct_col_o;
wire                      ct_gecerli_o;
wire                      ct_hazir_i = 1;
wire                      ct_blok_son_o;

huffman_decoder uut (
    .clk_i         ( clk_i ),
    .rstn_i        ( rstn_i ),
    .m_veri_i      ( m_veri_i ),
    .m_gecerli_i   ( m_gecerli_i ),
    .m_hazir_o     ( m_hazir_o ),
    .nd_run_o      ( nd_run_o ),
    .nd_data_o     ( nd_data_o ),
    .nd_gecerli_o  ( nd_gecerli_o ),
    .nd_hazir_i    ( nd_hazir_i ),
    .nd_blk_son_o  ( nd_blk_son_o )
);

zigzag_normalizer zn (
    .clk_i         ( clk_i ),
    .rstn_i        ( rstn_i ),
    .blok_son_i    ( nd_blk_son_o ),
    .hd_run_i      ( nd_run_o ),
    .hd_veri_i     ( nd_data_o ),
    .hd_gecerli_i  ( nd_gecerli_o ),
    .hd_hazir_o    ( nd_hazir_i ),
    .ct_veri_o     ( ct_veri_o ),
    .ct_row_o      ( ct_row_o ),
    .ct_col_o      ( ct_col_o ),
    .ct_gecerli_o  ( ct_gecerli_o ),
    .ct_blok_son_o ( ct_blok_son_o ),
    .ct_hazir_i    ( dq_zig_veri_hazir_w )
);

wire                      dq_zig_veri_hazir_w;
wire  [`Q_BIT-1:0]        dq_idct_veri_w;
wire  [`BLOCK_BIT-1:0]    dq_idct_veri_row_w;
wire  [`BLOCK_BIT-1:0]    dq_idct_veri_col_w;
wire                      dq_idct_veri_gecerli_w;
wire                      dq_idct_blok_son_w;
wire ict_dq_hazir_w;

dequantizer dq (
    .clk_i               ( clk_i ),
    .rstn_i              ( rstn_i ),
    .zig_veri_i          ( ct_veri_o ),
    .zig_veri_row_i      ( ct_row_o ),
    .zig_veri_col_i      ( ct_col_o ),
    .zig_veri_gecerli_i  ( ct_gecerli_o ),
    .zig_blok_son_i      ( ct_blok_son_o ),
    .zig_veri_hazir_o    ( dq_zig_veri_hazir_w ),
    .idct_veri_o         ( dq_idct_veri_w ),
    .idct_veri_row_o     ( dq_idct_veri_row_w ),
    .idct_veri_col_o     ( dq_idct_veri_col_w ),
    .idct_veri_gecerli_o ( dq_idct_veri_gecerli_w ),
    .idct_blok_son_o     ( dq_idct_blok_son_w ),
    .idct_veri_hazir_i   ( ict_dq_hazir_w )
);

wire                      ict_dq_hazir_w;
wire  [`PIXEL_BIT-1:0]    ict_gd_veri_w;
wire  [`BLOCK_BIT-1:0]    ict_gd_row_w;
wire  [`BLOCK_BIT-1:0]    ict_gd_col_w;
wire                      ict_gd_gecerli_w;
wire                      ict_gd_blok_son_w;

icosine_transformer ict (
    .clk_i          ( clk_i ),
    .rstn_i         ( rstn_i ),
    .dq_veri_i      ( dq_idct_veri_w ),
    .dq_row_i       ( dq_idct_veri_row_w ),
    .dq_col_i       ( dq_idct_veri_col_w ),
    .dq_gecerli_i   ( dq_idct_veri_gecerli_w ),
    .dq_blok_son_i  ( dq_idct_blok_son_w ),
    .dq_hazir_o     ( ict_dq_hazir_w ),
    .gd_veri_o      ( ict_gd_veri_w ),
    .gd_row_o       ( ict_gd_row_w ),
    .gd_col_o       ( ict_gd_col_w ),
    .gd_gecerli_o   ( ict_gd_gecerli_w ),
    .gd_blok_son_o  ( ict_gd_blok_son_w ),
    .gd_hazir_i     ( idct_hazir_w )
);

wire idct_hazir_w;
wire[7:0] coz_veri_o;
wire coz_gecerli_o;
wire coz_hazir_i =1;

decode_normalizer denorm (
    .clk_i           ( clk_i ),
    .rstn_i          ( rstn_i ),
    .idct_veri_i     ( ict_gd_veri_w ),
    .idct_row_i      ( ict_gd_row_w ),
    .idct_col_i      ( ict_gd_col_w ),
    .idct_gecerli_i  ( ict_gd_gecerli_w ),
    .idct_blok_son_i ( ict_gd_blok_son_w ),
    .idct_hazir_o    ( idct_hazir_w ),
    .dn_veri_o       ( coz_veri_o ),
    .dn_gecerli_o    ( coz_gecerli_o ),
    .dn_hazir_i      ( coz_hazir_i )
);

always begin
    clk_i = 1'b1;
    #5;
    clk_i = 1'b0;
    #5;
end

localparam TEST_LEN = 144;
localparam BYTE_LEN = TEST_LEN/8;
reg [TEST_LEN-1:0] temp_deger;
reg [7:0] bytes [0:BYTE_LEN-1];

integer step;

integer i;
initial begin
    dc_ready_i = 1;
    step = 0;
    temp_deger = 144'b101101000111111101110111111111110001111100110101011010001111111011101111111111100011111001101010110100011111110111011111111111000111110011010000;
    //temp_deger = 8072'b11100010000101011000101011110000011110100101001010110110000110111001110011110011111011110100111010001011100001110001100100111100010100111001110100110000110110001110001010010000001000011010100101000000001110000000001110000011010011010010000001110111110011111101011010011010110100001000001000001110000011110011111111001110101000010010000010000011100000111101010001010011100000110111101010001100110100000001010000011010100110111000001100010110001110111000111010110100100010101001100110101001010101100011001010100011001011000000100000000110101000101001010000011100110101000010011110000011010011111000100011100001101110100101010010001100100001000001101001010000110000000010111110111101001100011011001001110000011010100101100010001110000010001110011110001010001001010100110010110001101001001000110001111100111001010111000000001000001000101010001101110001101101011011000001101001010000001110011100110100111001110001110000000011010100011011110101000111110111101001110000111010110100111111011011110001100110100110111101111010001100011101011010011001100011111001101010000011010000101000110011010100100001111110010100011110111101010001111000110010011010101100110110111010111100110001100100011110101110011010010110011001111100101100111011011111100111010101010011101010011100010101001010110100001001111001110001110011111011010100110000000010100111111011011110001111011010100111011000000001110001110011110010001010100100100011100101000000110010000001110000011100011100000100110100100110111001101100100101101100111001110011010010000010010100011001110000010001111110010101010010001010000101011000000000111000111110101101001101100100100011010011100011000001111110101111011010101000000110010000001010011110000011100100010100101010100000000100011000110011010011100001110000001100111101011010010100001110010100111010000010100111101100110111100110000111100100100111100111101101110110101001101100100111001010111100100011100100011101111010100001011001011110011010010110001100011100110101011110011001000001001001000000000111010100000011001000001110110100111111110100101010100101001001111101111010100111101000001100101001111101001010011111000110001100000000110101001100111001110111001010001110001110011010100001100100010011011010110111000101010001000100111011100001100111101111010000000011010100100001111001100011001101010001000100011100010100110100100010100000000011100110101001010110111000000000000101010001111101111010000001110111101001101110001110011100110100100110001100110101001000101000110000001010010011000001001001110011010000000000000000011100011101110011010101101011001000010100000011011011110101000101010101100110001001001000001101001100010100000000011001001101010111010111010010000001101100011011000111111111010010101010110011010001000111100111000001110010011110110111101111010011000000010010001110001110111101001110001110001100100000100000111000001111011110100111111000010100111100100001100001010011100101011000011101000010101000000111110100101001101001000000111001111000101001010001001000110010111000111000110010001010100101001101110000101011000011111001100101001001001111010011001101001100011001010100011011100101010000011111101001010100010011001011101101001110010001110010001111111001010100101000111000111011010100000011100100111000101010010001011100101011110100001111000111101000011010011110111001010101100101111010100011001110001111010010100110001100000000110001001110001110100111101011010100011000000110000011110110101001111000100101001010011001000000111010001101110101000101001101110001101110011111001111010110101001001000100101110000100011000011101111010011101101101110110011000111111010110101011000100100100000001000010000011110101111011010101010110100100000110001100010101000100110010111100000111000000101001101000111010010101001011000110001100101010010001111011010100110100101011100100010101000110110000110001010010001010001111100110101001111011100110100110011101111010010110100110111000101000010100011100110101001110100100010110111000011001001001000000000110000010011010100011011111000111011000000100010100110101010001100001101111101001010011111101111001000000011011110101001101001000000101111110010100110101000110110000110001010011110101100101000111011101011100110101001000111011101010111010111000000011011000101010000101100101001001111010100111100110100100000110010000011110100110011010011111100100000100011111011101110001010011100100010111001111001000110011110001110101101001010010101110011110110101001111100011010100000100000100000110100100011101001100011111011101000110011010010000001100010001110101000001101001101001110000010011110000011010011101101101001110001100011101101010011101000111000111100101101010101100110010101000000101010000000111000000001111101001111011110101010100011001000010101011010100111000001111101101011011000111001001000001111011010100001100101110111000100111000000110001010100011110000010010011010101100110110111100010001011000011001111011110100010011101011101100100100000011001010110110010001100011100100010100100010100100101111100011111101001110001010101110010010110010011111101110110101000000110000011001001100011000110010001110110000101010101010110010100011000001000000111010010101000110000101110001100100011110101101010001111011011100011100000100011100110100101000001110001110001010011110101000111110010100110101000010111000110001010011010100000110010110101001010111111010110100100010000011001011010100101011010100110100110100101000101001111011010010000100100011000111010000011000101010001100100100100110100111100000011000010100100111110100110001010011010100000001011000100100111101110011110100101001111001000110000001100011101010010001110110101000110110001010000101110010110001111001001111011010101010111000111010110100111011101010001100111110100101000010100100100011111010010101001000001100101101100000100000101011010010100100000100111110100111111000010100101010000100101000011110101001111111000010100111100011100100110100111101010101001110011100100010100101011101011100011111111111010110101010001100101001110001100100000100111110111101001101110110111000101010011101001100000101011110010001010011101000110000000101011000111110111101001000001100101100010010101111111010010100111101011000011101111011000000011101110011010011001001101000011100001010110110001110101010110100110101010011101110010100000000100111111001100001110111101001110010110001000100111110100110001010100110001001000100001000111110100111001010110101000010001111100111000110110100011101010010011100111001111101011010100101010010000100110001110001001101001000011100111100000011100011111010110100100100011110010110001111111000011000101001011001000100001010100010101010110001001110010010110111001101010011010111001100010111010001101110001100111000111001101010000000000000011100111001101010010001000001100101010011010100000100101000111001101001100010011100011100110100100011011100110100111010001100011000000001001101001101001111010110100100110001010000011010001100110100011101100011010011110111111001000011000111101100000011010010001000001100000100011110101001000110011010011100000001101101110010000001111101111010100110001101100100000010100100001010111001000111000000111001101001101000111101001010011101101101101001110010000011000001000110010001110001010100110011001000000001110100111001000101001101001000110011110110101001010100111110010101101110011110100101010011001100000000000001110101000001111101000010001010011010111011011001111010010100101100011011011000111000101001110110110011001000110010001110001111011010100001100101110001110010001010010001010000000110001111010110101001010101000000010101110001100000111111100011100010101001011101111000110110111011101100011100111101111010100010100100011000001110110000011011111110000111000101001100010110000101100110011011100000011101011010100100110011101101011100101000001110100010111101001010100011100110110111010010001110000010000001110000000001100010100110110000101011110011100000000111000110011010101111010111001111111011110110110110010011000001110001101101111010100000011101111111011110101010111010111111101110110111111101100011010100100100101001000110110111100010101010101110110100011001111001000101010010100111001001010000;
    for (i = 0; i < BYTE_LEN; i = i + 1) begin
        bytes[i] = temp_deger[TEST_LEN - 1 - 8 * i -: 8];
    end
    rstn_i = 1'b0;
    m_gecerli_i = 0;
    repeat(20) @(posedge clk_i);
    rstn_i = 1'b1;

    for (i = 0; i < BYTE_LEN;) begin
        m_veri_i = bytes[i];
        m_gecerli_i = 1;
        @(posedge clk_i); #2;
        if (m_gecerli_i && m_hazir_o) begin
            i = i + 1;
        end
    end
    m_gecerli_i = 1'b0;
end

endmodule